module Registradores(r0enable, bus, clock, r0out);
	input r0enable;
	input [15:0]bus;
	input clock;
	output [15:0]r0out;



endmodule